`timescale 1ns / 1ps
module instmem(instr_addr,instruction);
input [31:0] instr_addr;
output [31:0] instruction;
reg[31:0] instruction;
reg [7:0] ram [90:0];
initial
  begin
    ram[0]  = 8'b00010011;
ram[1]  = 8'b00000000;
ram[2]  = 8'b10100000;
ram[3]  = 8'b00000000;

ram[4]  = 8'b10010011;
ram[5]  = 8'b00000101;
ram[6]  = 8'b01010000;
ram[7]  = 8'b00000000;

ram[8]  = 8'b00010011;
ram[9]  = 8'b00000000;
ram[10] = 8'b11110000;
ram[11] = 8'b00000000;

ram[12] = 8'b10110011;
ram[13] = 8'b10000001;
ram[14] = 8'b00100000;
ram[15] = 8'b00000000;

ram[16] = 8'b00110011;
ram[17] = 8'b10100010;
ram[18] = 8'b00110001;
ram[19] = 8'b00000000;

ram[20] = 8'b00110011;
ram[21] = 8'b10110010;
ram[22] = 8'b00110001;
ram[23] = 8'b00000000;

ram[24] = 8'b00110011;
ram[25] = 8'b10110011;
ram[26] = 8'b01100010;
ram[27] = 8'b00000000;

ram[28] = 8'b10110011;
ram[29] = 8'b10110011;
ram[30] = 8'b00100011;
ram[31] = 8'b00000000;

ram[32] = 8'b10110011;
ram[33] = 8'b11000011;
ram[34] = 8'b00010011;
ram[35] = 8'b00000000;

ram[36] = 8'b00100011;
ram[37] = 8'b00100000;
ram[38] = 8'b01000001;
ram[39] = 8'b00000000;

ram[40] = 8'b10100011;
ram[41] = 8'b00100000;
ram[42] = 8'b01010001;
ram[43] = 8'b00000000;

ram[44] = 8'b10000011;
ram[45] = 8'b00100010;
ram[46] = 8'b00000001;
ram[47] = 8'b00000000;

ram[48] = 8'b00000011;
ram[49] = 8'b00100011;
ram[50] = 8'b01000001;
ram[51] = 8'b00000000;

ram[52] = 8'b00110011;
ram[53] = 8'b01100011;
ram[54] = 8'b10110010;
ram[55] = 8'b00000000;

ram[56] = 8'b11100011;
ram[57] = 8'b00011100;
ram[58] = 8'b00100010;
ram[59] = 8'b11111110;

ram[60] = 8'b10010011;
ram[61] = 8'b00000110;
ram[62] = 8'b11111111;
ram[63] = 8'b00000000;

ram[64] = 8'b00110011;
ram[65] = 8'b01100011;
ram[66] = 8'b10100011;
ram[67] = 8'b01000000;

ram[68] = 8'b10110011;
ram[69] = 8'b11100011;
ram[70] = 8'b00110011;
ram[71] = 8'b00000000;

  end
    always @(instr_addr)
instruction = {ram[instr_addr+3],ram[instr_addr+2],ram[instr_addr+1],ram[instr_addr]};
endmodule
